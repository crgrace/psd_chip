// File Name: regfile_assign.sv
// Engineer:  Carl Grace (crgrace@lbl.gov)
// Description:  Code used in regfile.sv for assignment
//          
///////////////////////////////////////////////////////////////////

 
config_bits[CHANNEL_DISABLE] <= 8'h00;
config_bits[BUFF_REF0] <= 8'h00;
config_bits[BUFF_REF1] <= 8'h00;
config_bits[BUFF_REF2] <= 8'h00;
config_bits[BUFF_REF3] <= 8'h00;
config_bits[BUFF_REF4] <= 8'h00;
config_bits[D2S_REF0] <= 8'h00;
config_bits[D2S_REF1] <= 8'h00;
config_bits[D2S_REF2] <= 8'h00;
config_bits[D2S_REF3] <= 8'h00;
config_bits[THRESH_SOUT_GLOBAL] <= 8'h00;
config_bits[THRESH_SOUT_FINE0] <= 8'h00;
config_bits[THRESH_SOUT_FINE1] <= 8'h00;
config_bits[THRESH_SOUT_FINE2] <= 8'h00;
config_bits[THRESH_SOUT_FINE3] <= 8'h00;
config_bits[THRESH_FOUT_GLOBAL] <= 8'h00;
config_bits[THRESH_FOUT_FINE0] <= 8'h00;
config_bits[THRESH_FOUT_FINE1] <= 8'h00;
config_bits[THRESH_FOUT_FINE2] <= 8'h00;
config_bits[THRESH_FOUT_FINE3] <= 8'h00;
config_bits[IBIAS_TOTAL_INT] <= 8'h00;
config_bits[IBIAS_PARTIAL_INT] <= 8'h00;
config_bits[IBIAS_DISC] <= 8'h00;
config_bits[IBIAS_DISC_OUT] <= 8'h00;
config_bits[IBIAS_FOUT_WIDTH] <= 8'h00;
config_bits[IBIAS_LVDS] <= 8'h00;
config_bits[TUNABLE_RES_TOTAL_INT] <= 8'h00;
config_bits[TUNABLE_RES_SUBTR_GAIN] <= 8'h00;
config_bits[SEL_WIDTH] <= 8'h00;
config_bits[IMONITOR] <= 8'h00;
config_bits[VMONITOR] <= 8'h00;


